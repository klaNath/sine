						
module	diff_rom	(
    input	wire	[8:0]	inadrs, 	
    output	wire	[15:0]	outdiff);		
						
	assign	outdiff = sin_rom(inadrs);				
						
	function	[15:0]	sin_rom;			
						
		input	[8:0]	adrs;		
		begin				
		case	(adrs)			
		9'D0	:	sin_rom =	201	;
		9'D1	:	sin_rom =	201	;
		9'D2	:	sin_rom =	202	;
		9'D3	:	sin_rom =	201	;
		9'D4	:	sin_rom =	202	;
		9'D5	:	sin_rom =	201	;
		9'D6	:	sin_rom =	202	;
		9'D7	:	sin_rom =	201	;
		9'D8	:	sin_rom =	201	;
		9'D9	:	sin_rom =	202	;
		9'D10	:	sin_rom =	201	;
		9'D11	:	sin_rom =	201	;
		9'D12	:	sin_rom =	202	;
		9'D13	:	sin_rom =	201	;
		9'D14	:	sin_rom =	201	;
		9'D15	:	sin_rom =	201	;
		9'D16	:	sin_rom =	202	;
		9'D17	:	sin_rom =	201	;
		9'D18	:	sin_rom =	201	;
		9'D19	:	sin_rom =	201	;
		9'D20	:	sin_rom =	201	;
		9'D21	:	sin_rom =	201	;
		9'D22	:	sin_rom =	201	;
		9'D23	:	sin_rom =	201	;
		9'D24	:	sin_rom =	201	;
		9'D25	:	sin_rom =	201	;
		9'D26	:	sin_rom =	201	;
		9'D27	:	sin_rom =	200	;
		9'D28	:	sin_rom =	201	;
		9'D29	:	sin_rom =	201	;
		9'D30	:	sin_rom =	200	;
		9'D31	:	sin_rom =	201	;
		9'D32	:	sin_rom =	200	;
		9'D33	:	sin_rom =	201	;
		9'D34	:	sin_rom =	200	;
		9'D35	:	sin_rom =	200	;
		9'D36	:	sin_rom =	200	;
		9'D37	:	sin_rom =	200	;
		9'D38	:	sin_rom =	200	;
		9'D39	:	sin_rom =	200	;
		9'D40	:	sin_rom =	200	;
		9'D41	:	sin_rom =	200	;
		9'D42	:	sin_rom =	200	;
		9'D43	:	sin_rom =	200	;
		9'D44	:	sin_rom =	199	;
		9'D45	:	sin_rom =	200	;
		9'D46	:	sin_rom =	199	;
		9'D47	:	sin_rom =	199	;
		9'D48	:	sin_rom =	200	;
		9'D49	:	sin_rom =	199	;
		9'D50	:	sin_rom =	199	;
		9'D51	:	sin_rom =	199	;
		9'D52	:	sin_rom =	198	;
		9'D53	:	sin_rom =	199	;
		9'D54	:	sin_rom =	199	;
		9'D55	:	sin_rom =	198	;
		9'D56	:	sin_rom =	199	;
		9'D57	:	sin_rom =	198	;
		9'D58	:	sin_rom =	198	;
		9'D59	:	sin_rom =	198	;
		9'D60	:	sin_rom =	198	;
		9'D61	:	sin_rom =	198	;
		9'D62	:	sin_rom =	198	;
		9'D63	:	sin_rom =	198	;
		9'D64	:	sin_rom =	197	;
		9'D65	:	sin_rom =	198	;
		9'D66	:	sin_rom =	197	;
		9'D67	:	sin_rom =	197	;
		9'D68	:	sin_rom =	197	;
		9'D69	:	sin_rom =	197	;
		9'D70	:	sin_rom =	197	;
		9'D71	:	sin_rom =	196	;
		9'D72	:	sin_rom =	197	;
		9'D73	:	sin_rom =	196	;
		9'D74	:	sin_rom =	196	;
		9'D75	:	sin_rom =	196	;
		9'D76	:	sin_rom =	196	;
		9'D77	:	sin_rom =	196	;
		9'D78	:	sin_rom =	196	;
		9'D79	:	sin_rom =	195	;
		9'D80	:	sin_rom =	195	;
		9'D81	:	sin_rom =	195	;
		9'D82	:	sin_rom =	195	;
		9'D83	:	sin_rom =	195	;
		9'D84	:	sin_rom =	195	;
		9'D85	:	sin_rom =	195	;
		9'D86	:	sin_rom =	194	;
		9'D87	:	sin_rom =	194	;
		9'D88	:	sin_rom =	194	;
		9'D89	:	sin_rom =	194	;
		9'D90	:	sin_rom =	194	;
		9'D91	:	sin_rom =	193	;
		9'D92	:	sin_rom =	194	;
		9'D93	:	sin_rom =	193	;
		9'D94	:	sin_rom =	193	;
		9'D95	:	sin_rom =	193	;
		9'D96	:	sin_rom =	192	;
		9'D97	:	sin_rom =	193	;
		9'D98	:	sin_rom =	192	;
		9'D99	:	sin_rom =	192	;
		9'D100	:	sin_rom =	192	;
		9'D101	:	sin_rom =	192	;
		9'D102	:	sin_rom =	191	;
		9'D103	:	sin_rom =	192	;
		9'D104	:	sin_rom =	191	;
		9'D105	:	sin_rom =	191	;
		9'D106	:	sin_rom =	191	;
		9'D107	:	sin_rom =	190	;
		9'D108	:	sin_rom =	191	;
		9'D109	:	sin_rom =	190	;
		9'D110	:	sin_rom =	190	;
		9'D111	:	sin_rom =	189	;
		9'D112	:	sin_rom =	190	;
		9'D113	:	sin_rom =	189	;
		9'D114	:	sin_rom =	189	;
		9'D115	:	sin_rom =	189	;
		9'D116	:	sin_rom =	189	;
		9'D117	:	sin_rom =	188	;
		9'D118	:	sin_rom =	189	;
		9'D119	:	sin_rom =	188	;
		9'D120	:	sin_rom =	187	;
		9'D121	:	sin_rom =	188	;
		9'D122	:	sin_rom =	187	;
		9'D123	:	sin_rom =	187	;
		9'D124	:	sin_rom =	187	;
		9'D125	:	sin_rom =	187	;
		9'D126	:	sin_rom =	186	;
		9'D127	:	sin_rom =	187	;
		9'D128	:	sin_rom =	186	;
		9'D129	:	sin_rom =	185	;
		9'D130	:	sin_rom =	186	;
		9'D131	:	sin_rom =	185	;
		9'D132	:	sin_rom =	185	;
		9'D133	:	sin_rom =	185	;
		9'D134	:	sin_rom =	184	;
		9'D135	:	sin_rom =	184	;
		9'D136	:	sin_rom =	184	;
		9'D137	:	sin_rom =	184	;
		9'D138	:	sin_rom =	183	;
		9'D139	:	sin_rom =	184	;
		9'D140	:	sin_rom =	183	;
		9'D141	:	sin_rom =	182	;
		9'D142	:	sin_rom =	183	;
		9'D143	:	sin_rom =	182	;
		9'D144	:	sin_rom =	182	;
		9'D145	:	sin_rom =	182	;
		9'D146	:	sin_rom =	181	;
		9'D147	:	sin_rom =	181	;
		9'D148	:	sin_rom =	181	;
		9'D149	:	sin_rom =	180	;
		9'D150	:	sin_rom =	181	;
		9'D151	:	sin_rom =	180	;
		9'D152	:	sin_rom =	179	;
		9'D153	:	sin_rom =	180	;
		9'D154	:	sin_rom =	179	;
		9'D155	:	sin_rom =	179	;
		9'D156	:	sin_rom =	178	;
		9'D157	:	sin_rom =	179	;
		9'D158	:	sin_rom =	178	;
		9'D159	:	sin_rom =	177	;
		9'D160	:	sin_rom =	178	;
		9'D161	:	sin_rom =	177	;
		9'D162	:	sin_rom =	177	;
		9'D163	:	sin_rom =	176	;
		9'D164	:	sin_rom =	177	;
		9'D165	:	sin_rom =	176	;
		9'D166	:	sin_rom =	175	;
		9'D167	:	sin_rom =	176	;
		9'D168	:	sin_rom =	175	;
		9'D169	:	sin_rom =	174	;
		9'D170	:	sin_rom =	175	;
		9'D171	:	sin_rom =	174	;
		9'D172	:	sin_rom =	174	;
		9'D173	:	sin_rom =	173	;
		9'D174	:	sin_rom =	173	;
		9'D175	:	sin_rom =	173	;
		9'D176	:	sin_rom =	173	;
		9'D177	:	sin_rom =	172	;
		9'D178	:	sin_rom =	172	;
		9'D179	:	sin_rom =	171	;
		9'D180	:	sin_rom =	172	;
		9'D181	:	sin_rom =	170	;
		9'D182	:	sin_rom =	171	;
		9'D183	:	sin_rom =	170	;
		9'D184	:	sin_rom =	170	;
		9'D185	:	sin_rom =	170	;
		9'D186	:	sin_rom =	169	;
		9'D187	:	sin_rom =	169	;
		9'D188	:	sin_rom =	168	;
		9'D189	:	sin_rom =	169	;
		9'D190	:	sin_rom =	168	;
		9'D191	:	sin_rom =	167	;
		9'D192	:	sin_rom =	167	;
		9'D193	:	sin_rom =	167	;
		9'D194	:	sin_rom =	167	;
		9'D195	:	sin_rom =	166	;
		9'D196	:	sin_rom =	166	;
		9'D197	:	sin_rom =	165	;
		9'D198	:	sin_rom =	165	;
		9'D199	:	sin_rom =	165	;
		9'D200	:	sin_rom =	164	;
		9'D201	:	sin_rom =	164	;
		9'D202	:	sin_rom =	164	;
		9'D203	:	sin_rom =	163	;
		9'D204	:	sin_rom =	163	;
		9'D205	:	sin_rom =	163	;
		9'D206	:	sin_rom =	162	;
		9'D207	:	sin_rom =	162	;
		9'D208	:	sin_rom =	161	;
		9'D209	:	sin_rom =	162	;
		9'D210	:	sin_rom =	160	;
		9'D211	:	sin_rom =	161	;
		9'D212	:	sin_rom =	160	;
		9'D213	:	sin_rom =	159	;
		9'D214	:	sin_rom =	159	;
		9'D215	:	sin_rom =	159	;
		9'D216	:	sin_rom =	159	;
		9'D217	:	sin_rom =	158	;
		9'D218	:	sin_rom =	158	;
		9'D219	:	sin_rom =	157	;
		9'D220	:	sin_rom =	157	;
		9'D221	:	sin_rom =	156	;
		9'D222	:	sin_rom =	156	;
		9'D223	:	sin_rom =	156	;
		9'D224	:	sin_rom =	156	;
		9'D225	:	sin_rom =	155	;
		9'D226	:	sin_rom =	154	;
		9'D227	:	sin_rom =	154	;
		9'D228	:	sin_rom =	154	;
		9'D229	:	sin_rom =	153	;
		9'D230	:	sin_rom =	153	;
		9'D231	:	sin_rom =	153	;
		9'D232	:	sin_rom =	152	;
		9'D233	:	sin_rom =	152	;
		9'D234	:	sin_rom =	151	;
		9'D235	:	sin_rom =	151	;
		9'D236	:	sin_rom =	151	;
		9'D237	:	sin_rom =	150	;
		9'D238	:	sin_rom =	149	;
		9'D239	:	sin_rom =	150	;
		9'D240	:	sin_rom =	149	;
		9'D241	:	sin_rom =	148	;
		9'D242	:	sin_rom =	148	;
		9'D243	:	sin_rom =	148	;
		9'D244	:	sin_rom =	147	;
		9'D245	:	sin_rom =	147	;
		9'D246	:	sin_rom =	146	;
		9'D247	:	sin_rom =	146	;
		9'D248	:	sin_rom =	145	;
		9'D249	:	sin_rom =	145	;
		9'D250	:	sin_rom =	145	;
		9'D251	:	sin_rom =	144	;
		9'D252	:	sin_rom =	144	;
		9'D253	:	sin_rom =	143	;
		9'D254	:	sin_rom =	143	;
		9'D255	:	sin_rom =	143	;
		9'D256	:	sin_rom =	142	;
		9'D257	:	sin_rom =	141	;
		9'D258	:	sin_rom =	141	;
		9'D259	:	sin_rom =	141	;
		9'D260	:	sin_rom =	140	;
		9'D261	:	sin_rom =	140	;
		9'D262	:	sin_rom =	139	;
		9'D263	:	sin_rom =	139	;
		9'D264	:	sin_rom =	139	;
		9'D265	:	sin_rom =	138	;
		9'D266	:	sin_rom =	137	;
		9'D267	:	sin_rom =	137	;
		9'D268	:	sin_rom =	137	;
		9'D269	:	sin_rom =	136	;
		9'D270	:	sin_rom =	136	;
		9'D271	:	sin_rom =	135	;
		9'D272	:	sin_rom =	135	;
		9'D273	:	sin_rom =	134	;
		9'D274	:	sin_rom =	134	;
		9'D275	:	sin_rom =	134	;
		9'D276	:	sin_rom =	133	;
		9'D277	:	sin_rom =	132	;
		9'D278	:	sin_rom =	132	;
		9'D279	:	sin_rom =	132	;
		9'D280	:	sin_rom =	131	;
		9'D281	:	sin_rom =	131	;
		9'D282	:	sin_rom =	130	;
		9'D283	:	sin_rom =	129	;
		9'D284	:	sin_rom =	130	;
		9'D285	:	sin_rom =	128	;
		9'D286	:	sin_rom =	129	;
		9'D287	:	sin_rom =	127	;
		9'D288	:	sin_rom =	128	;
		9'D289	:	sin_rom =	126	;
		9'D290	:	sin_rom =	127	;
		9'D291	:	sin_rom =	126	;
		9'D292	:	sin_rom =	125	;
		9'D293	:	sin_rom =	125	;
		9'D294	:	sin_rom =	124	;
		9'D295	:	sin_rom =	124	;
		9'D296	:	sin_rom =	124	;
		9'D297	:	sin_rom =	122	;
		9'D298	:	sin_rom =	123	;
		9'D299	:	sin_rom =	122	;
		9'D300	:	sin_rom =	121	;
		9'D301	:	sin_rom =	121	;
		9'D302	:	sin_rom =	121	;
		9'D303	:	sin_rom =	120	;
		9'D304	:	sin_rom =	119	;
		9'D305	:	sin_rom =	119	;
		9'D306	:	sin_rom =	119	;
		9'D307	:	sin_rom =	118	;
		9'D308	:	sin_rom =	117	;
		9'D309	:	sin_rom =	117	;
		9'D310	:	sin_rom =	116	;
		9'D311	:	sin_rom =	116	;
		9'D312	:	sin_rom =	116	;
		9'D313	:	sin_rom =	115	;
		9'D314	:	sin_rom =	114	;
		9'D315	:	sin_rom =	114	;
		9'D316	:	sin_rom =	113	;
		9'D317	:	sin_rom =	113	;
		9'D318	:	sin_rom =	113	;
		9'D319	:	sin_rom =	112	;
		9'D320	:	sin_rom =	111	;
		9'D321	:	sin_rom =	111	;
		9'D322	:	sin_rom =	110	;
		9'D323	:	sin_rom =	110	;
		9'D324	:	sin_rom =	109	;
		9'D325	:	sin_rom =	109	;
		9'D326	:	sin_rom =	108	;
		9'D327	:	sin_rom =	108	;
		9'D328	:	sin_rom =	107	;
		9'D329	:	sin_rom =	107	;
		9'D330	:	sin_rom =	106	;
		9'D331	:	sin_rom =	105	;
		9'D332	:	sin_rom =	105	;
		9'D333	:	sin_rom =	105	;
		9'D334	:	sin_rom =	104	;
		9'D335	:	sin_rom =	103	;
		9'D336	:	sin_rom =	103	;
		9'D337	:	sin_rom =	103	;
		9'D338	:	sin_rom =	102	;
		9'D339	:	sin_rom =	101	;
		9'D340	:	sin_rom =	101	;
		9'D341	:	sin_rom =	100	;
		9'D342	:	sin_rom =	100	;
		9'D343	:	sin_rom =	99	;
		9'D344	:	sin_rom =	99	;
		9'D345	:	sin_rom =	98	;
		9'D346	:	sin_rom =	97	;
		9'D347	:	sin_rom =	98	;
		9'D348	:	sin_rom =	96	;
		9'D349	:	sin_rom =	96	;
		9'D350	:	sin_rom =	95	;
		9'D351	:	sin_rom =	95	;
		9'D352	:	sin_rom =	95	;
		9'D353	:	sin_rom =	93	;
		9'D354	:	sin_rom =	94	;
		9'D355	:	sin_rom =	92	;
		9'D356	:	sin_rom =	92	;
		9'D357	:	sin_rom =	92	;
		9'D358	:	sin_rom =	91	;
		9'D359	:	sin_rom =	90	;
		9'D360	:	sin_rom =	90	;
		9'D361	:	sin_rom =	90	;
		9'D362	:	sin_rom =	88	;
		9'D363	:	sin_rom =	89	;
		9'D364	:	sin_rom =	87	;
		9'D365	:	sin_rom =	88	;
		9'D366	:	sin_rom =	86	;
		9'D367	:	sin_rom =	86	;
		9'D368	:	sin_rom =	86	;
		9'D369	:	sin_rom =	84	;
		9'D370	:	sin_rom =	85	;
		9'D371	:	sin_rom =	84	;
		9'D372	:	sin_rom =	83	;
		9'D373	:	sin_rom =	82	;
		9'D374	:	sin_rom =	82	;
		9'D375	:	sin_rom =	82	;
		9'D376	:	sin_rom =	81	;
		9'D377	:	sin_rom =	80	;
		9'D378	:	sin_rom =	80	;
		9'D379	:	sin_rom =	79	;
		9'D380	:	sin_rom =	79	;
		9'D381	:	sin_rom =	78	;
		9'D382	:	sin_rom =	78	;
		9'D383	:	sin_rom =	77	;
		9'D384	:	sin_rom =	76	;
		9'D385	:	sin_rom =	76	;
		9'D386	:	sin_rom =	75	;
		9'D387	:	sin_rom =	75	;
		9'D388	:	sin_rom =	74	;
		9'D389	:	sin_rom =	73	;
		9'D390	:	sin_rom =	73	;
		9'D391	:	sin_rom =	72	;
		9'D392	:	sin_rom =	72	;
		9'D393	:	sin_rom =	71	;
		9'D394	:	sin_rom =	71	;
		9'D395	:	sin_rom =	70	;
		9'D396	:	sin_rom =	70	;
		9'D397	:	sin_rom =	68	;
		9'D398	:	sin_rom =	69	;
		9'D399	:	sin_rom =	67	;
		9'D400	:	sin_rom =	67	;
		9'D401	:	sin_rom =	67	;
		9'D402	:	sin_rom =	66	;
		9'D403	:	sin_rom =	65	;
		9'D404	:	sin_rom =	65	;
		9'D405	:	sin_rom =	64	;
		9'D406	:	sin_rom =	64	;
		9'D407	:	sin_rom =	63	;
		9'D408	:	sin_rom =	62	;
		9'D409	:	sin_rom =	62	;
		9'D410	:	sin_rom =	61	;
		9'D411	:	sin_rom =	61	;
		9'D412	:	sin_rom =	60	;
		9'D413	:	sin_rom =	60	;
		9'D414	:	sin_rom =	59	;
		9'D415	:	sin_rom =	58	;
		9'D416	:	sin_rom =	58	;
		9'D417	:	sin_rom =	57	;
		9'D418	:	sin_rom =	56	;
		9'D419	:	sin_rom =	56	;
		9'D420	:	sin_rom =	55	;
		9'D421	:	sin_rom =	55	;
		9'D422	:	sin_rom =	54	;
		9'D423	:	sin_rom =	54	;
		9'D424	:	sin_rom =	53	;
		9'D425	:	sin_rom =	52	;
		9'D426	:	sin_rom =	52	;
		9'D427	:	sin_rom =	51	;
		9'D428	:	sin_rom =	51	;
		9'D429	:	sin_rom =	49	;
		9'D430	:	sin_rom =	50	;
		9'D431	:	sin_rom =	49	;
		9'D432	:	sin_rom =	48	;
		9'D433	:	sin_rom =	47	;
		9'D434	:	sin_rom =	47	;
		9'D435	:	sin_rom =	47	;
		9'D436	:	sin_rom =	45	;
		9'D437	:	sin_rom =	45	;
		9'D438	:	sin_rom =	45	;
		9'D439	:	sin_rom =	44	;
		9'D440	:	sin_rom =	43	;
		9'D441	:	sin_rom =	43	;
		9'D442	:	sin_rom =	42	;
		9'D443	:	sin_rom =	41	;
		9'D444	:	sin_rom =	41	;
		9'D445	:	sin_rom =	41	;
		9'D446	:	sin_rom =	39	;
		9'D447	:	sin_rom =	39	;
		9'D448	:	sin_rom =	39	;
		9'D449	:	sin_rom =	38	;
		9'D450	:	sin_rom =	37	;
		9'D451	:	sin_rom =	37	;
		9'D452	:	sin_rom =	36	;
		9'D453	:	sin_rom =	35	;
		9'D454	:	sin_rom =	35	;
		9'D455	:	sin_rom =	34	;
		9'D456	:	sin_rom =	34	;
		9'D457	:	sin_rom =	33	;
		9'D458	:	sin_rom =	32	;
		9'D459	:	sin_rom =	32	;
		9'D460	:	sin_rom =	31	;
		9'D461	:	sin_rom =	30	;
		9'D462	:	sin_rom =	30	;
		9'D463	:	sin_rom =	30	;
		9'D464	:	sin_rom =	28	;
		9'D465	:	sin_rom =	28	;
		9'D466	:	sin_rom =	28	;
		9'D467	:	sin_rom =	27	;
		9'D468	:	sin_rom =	26	;
		9'D469	:	sin_rom =	26	;
		9'D470	:	sin_rom =	25	;
		9'D471	:	sin_rom =	24	;
		9'D472	:	sin_rom =	24	;
		9'D473	:	sin_rom =	23	;
		9'D474	:	sin_rom =	23	;
		9'D475	:	sin_rom =	22	;
		9'D476	:	sin_rom =	21	;
		9'D477	:	sin_rom =	21	;
		9'D478	:	sin_rom =	20	;
		9'D479	:	sin_rom =	19	;
		9'D480	:	sin_rom =	19	;
		9'D481	:	sin_rom =	18	;
		9'D482	:	sin_rom =	18	;
		9'D483	:	sin_rom =	17	;
		9'D484	:	sin_rom =	16	;
		9'D485	:	sin_rom =	16	;
		9'D486	:	sin_rom =	15	;
		9'D487	:	sin_rom =	15	;
		9'D488	:	sin_rom =	14	;
		9'D489	:	sin_rom =	13	;
		9'D490	:	sin_rom =	13	;
		9'D491	:	sin_rom =	12	;
		9'D492	:	sin_rom =	11	;
		9'D493	:	sin_rom =	11	;
		9'D494	:	sin_rom =	10	;
		9'D495	:	sin_rom =	10	;
		9'D496	:	sin_rom =	9	;
		9'D497	:	sin_rom =	8	;
		9'D498	:	sin_rom =	8	;
		9'D499	:	sin_rom =	7	;
		9'D500	:	sin_rom =	7	;
		9'D501	:	sin_rom =	5	;
		9'D502	:	sin_rom =	6	;
		9'D503	:	sin_rom =	4	;
		9'D504	:	sin_rom =	4	;
		9'D505	:	sin_rom =	4	;
		9'D506	:	sin_rom =	3	;
		9'D507	:	sin_rom =	2	;
		9'D508	:	sin_rom =	1	;
		9'D509	:	sin_rom =	1	;
		9'D510	:	sin_rom =	1	;
		9'D511	:	sin_rom =	0	;
		default	:	sin_rom =	0	;
		endcase				
	end					
endfunction						
endmodule						
						
