						
module	sin_rom	(
    input	wire	[8:0]	inadrs, 	
    output	wire	[15:0]	outsine);			
							
	assign	outsine = sin_rom(inadrs);				
						
	function	[15:0]	sin_rom;			
						
		input	[8:0]	adrs;		
		begin				
		case	(adrs)			
		9'D0	:	sin_rom =	0	;
		9'D1	:	sin_rom =	201	;
		9'D2	:	sin_rom =	402	;
		9'D3	:	sin_rom =	604	;
		9'D4	:	sin_rom =	805	;
		9'D5	:	sin_rom =	1007	;
		9'D6	:	sin_rom =	1208	;
		9'D7	:	sin_rom =	1410	;
		9'D8	:	sin_rom =	1611	;
		9'D9	:	sin_rom =	1812	;
		9'D10	:	sin_rom =	2014	;
		9'D11	:	sin_rom =	2215	;
		9'D12	:	sin_rom =	2416	;
		9'D13	:	sin_rom =	2618	;
		9'D14	:	sin_rom =	2819	;
		9'D15	:	sin_rom =	3020	;
		9'D16	:	sin_rom =	3221	;
		9'D17	:	sin_rom =	3423	;
		9'D18	:	sin_rom =	3624	;
		9'D19	:	sin_rom =	3825	;
		9'D20	:	sin_rom =	4026	;
		9'D21	:	sin_rom =	4227	;
		9'D22	:	sin_rom =	4428	;
		9'D23	:	sin_rom =	4629	;
		9'D24	:	sin_rom =	4830	;
		9'D25	:	sin_rom =	5031	;
		9'D26	:	sin_rom =	5232	;
		9'D27	:	sin_rom =	5433	;
		9'D28	:	sin_rom =	5633	;
		9'D29	:	sin_rom =	5834	;
		9'D30	:	sin_rom =	6035	;
		9'D31	:	sin_rom =	6235	;
		9'D32	:	sin_rom =	6436	;
		9'D33	:	sin_rom =	6636	;
		9'D34	:	sin_rom =	6837	;
		9'D35	:	sin_rom =	7037	;
		9'D36	:	sin_rom =	7237	;
		9'D37	:	sin_rom =	7437	;
		9'D38	:	sin_rom =	7637	;
		9'D39	:	sin_rom =	7837	;
		9'D40	:	sin_rom =	8037	;
		9'D41	:	sin_rom =	8237	;
		9'D42	:	sin_rom =	8437	;
		9'D43	:	sin_rom =	8637	;
		9'D44	:	sin_rom =	8837	;
		9'D45	:	sin_rom =	9036	;
		9'D46	:	sin_rom =	9236	;
		9'D47	:	sin_rom =	9435	;
		9'D48	:	sin_rom =	9634	;
		9'D49	:	sin_rom =	9834	;
		9'D50	:	sin_rom =	10033	;
		9'D51	:	sin_rom =	10232	;
		9'D52	:	sin_rom =	10431	;
		9'D53	:	sin_rom =	10629	;
		9'D54	:	sin_rom =	10828	;
		9'D55	:	sin_rom =	11027	;
		9'D56	:	sin_rom =	11225	;
		9'D57	:	sin_rom =	11424	;
		9'D58	:	sin_rom =	11622	;
		9'D59	:	sin_rom =	11820	;
		9'D60	:	sin_rom =	12018	;
		9'D61	:	sin_rom =	12216	;
		9'D62	:	sin_rom =	12414	;
		9'D63	:	sin_rom =	12612	;
		9'D64	:	sin_rom =	12810	;
		9'D65	:	sin_rom =	13007	;
		9'D66	:	sin_rom =	13205	;
		9'D67	:	sin_rom =	13402	;
		9'D68	:	sin_rom =	13599	;
		9'D69	:	sin_rom =	13796	;
		9'D70	:	sin_rom =	13993	;
		9'D71	:	sin_rom =	14190	;
		9'D72	:	sin_rom =	14386	;
		9'D73	:	sin_rom =	14583	;
		9'D74	:	sin_rom =	14779	;
		9'D75	:	sin_rom =	14975	;
		9'D76	:	sin_rom =	15171	;
		9'D77	:	sin_rom =	15367	;
		9'D78	:	sin_rom =	15563	;
		9'D79	:	sin_rom =	15759	;
		9'D80	:	sin_rom =	15954	;
		9'D81	:	sin_rom =	16149	;
		9'D82	:	sin_rom =	16344	;
		9'D83	:	sin_rom =	16539	;
		9'D84	:	sin_rom =	16734	;
		9'D85	:	sin_rom =	16929	;
		9'D86	:	sin_rom =	17124	;
		9'D87	:	sin_rom =	17318	;
		9'D88	:	sin_rom =	17512	;
		9'D89	:	sin_rom =	17706	;
		9'D90	:	sin_rom =	17900	;
		9'D91	:	sin_rom =	18094	;
		9'D92	:	sin_rom =	18287	;
		9'D93	:	sin_rom =	18481	;
		9'D94	:	sin_rom =	18674	;
		9'D95	:	sin_rom =	18867	;
		9'D96	:	sin_rom =	19060	;
		9'D97	:	sin_rom =	19252	;
		9'D98	:	sin_rom =	19445	;
		9'D99	:	sin_rom =	19637	;
		9'D100	:	sin_rom =	19829	;
		9'D101	:	sin_rom =	20021	;
		9'D102	:	sin_rom =	20213	;
		9'D103	:	sin_rom =	20404	;
		9'D104	:	sin_rom =	20596	;
		9'D105	:	sin_rom =	20787	;
		9'D106	:	sin_rom =	20978	;
		9'D107	:	sin_rom =	21169	;
		9'D108	:	sin_rom =	21359	;
		9'D109	:	sin_rom =	21550	;
		9'D110	:	sin_rom =	21740	;
		9'D111	:	sin_rom =	21930	;
		9'D112	:	sin_rom =	22119	;
		9'D113	:	sin_rom =	22309	;
		9'D114	:	sin_rom =	22498	;
		9'D115	:	sin_rom =	22687	;
		9'D116	:	sin_rom =	22876	;
		9'D117	:	sin_rom =	23065	;
		9'D118	:	sin_rom =	23253	;
		9'D119	:	sin_rom =	23442	;
		9'D120	:	sin_rom =	23630	;
		9'D121	:	sin_rom =	23817	;
		9'D122	:	sin_rom =	24005	;
		9'D123	:	sin_rom =	24192	;
		9'D124	:	sin_rom =	24379	;
		9'D125	:	sin_rom =	24566	;
		9'D126	:	sin_rom =	24753	;
		9'D127	:	sin_rom =	24939	;
		9'D128	:	sin_rom =	25126	;
		9'D129	:	sin_rom =	25312	;
		9'D130	:	sin_rom =	25497	;
		9'D131	:	sin_rom =	25683	;
		9'D132	:	sin_rom =	25868	;
		9'D133	:	sin_rom =	26053	;
		9'D134	:	sin_rom =	26238	;
		9'D135	:	sin_rom =	26422	;
		9'D136	:	sin_rom =	26606	;
		9'D137	:	sin_rom =	26790	;
		9'D138	:	sin_rom =	26974	;
		9'D139	:	sin_rom =	27157	;
		9'D140	:	sin_rom =	27341	;
		9'D141	:	sin_rom =	27524	;
		9'D142	:	sin_rom =	27706	;
		9'D143	:	sin_rom =	27889	;
		9'D144	:	sin_rom =	28071	;
		9'D145	:	sin_rom =	28253	;
		9'D146	:	sin_rom =	28435	;
		9'D147	:	sin_rom =	28616	;
		9'D148	:	sin_rom =	28797	;
		9'D149	:	sin_rom =	28978	;
		9'D150	:	sin_rom =	29158	;
		9'D151	:	sin_rom =	29339	;
		9'D152	:	sin_rom =	29519	;
		9'D153	:	sin_rom =	29698	;
		9'D154	:	sin_rom =	29878	;
		9'D155	:	sin_rom =	30057	;
		9'D156	:	sin_rom =	30236	;
		9'D157	:	sin_rom =	30414	;
		9'D158	:	sin_rom =	30593	;
		9'D159	:	sin_rom =	30771	;
		9'D160	:	sin_rom =	30948	;
		9'D161	:	sin_rom =	31126	;
		9'D162	:	sin_rom =	31303	;
		9'D163	:	sin_rom =	31480	;
		9'D164	:	sin_rom =	31656	;
		9'D165	:	sin_rom =	31833	;
		9'D166	:	sin_rom =	32009	;
		9'D167	:	sin_rom =	32184	;
		9'D168	:	sin_rom =	32360	;
		9'D169	:	sin_rom =	32535	;
		9'D170	:	sin_rom =	32709	;
		9'D171	:	sin_rom =	32884	;
		9'D172	:	sin_rom =	33058	;
		9'D173	:	sin_rom =	33232	;
		9'D174	:	sin_rom =	33405	;
		9'D175	:	sin_rom =	33578	;
		9'D176	:	sin_rom =	33751	;
		9'D177	:	sin_rom =	33924	;
		9'D178	:	sin_rom =	34096	;
		9'D179	:	sin_rom =	34268	;
		9'D180	:	sin_rom =	34439	;
		9'D181	:	sin_rom =	34611	;
		9'D182	:	sin_rom =	34781	;
		9'D183	:	sin_rom =	34952	;
		9'D184	:	sin_rom =	35122	;
		9'D185	:	sin_rom =	35292	;
		9'D186	:	sin_rom =	35462	;
		9'D187	:	sin_rom =	35631	;
		9'D188	:	sin_rom =	35800	;
		9'D189	:	sin_rom =	35968	;
		9'D190	:	sin_rom =	36137	;
		9'D191	:	sin_rom =	36305	;
		9'D192	:	sin_rom =	36472	;
		9'D193	:	sin_rom =	36639	;
		9'D194	:	sin_rom =	36806	;
		9'D195	:	sin_rom =	36973	;
		9'D196	:	sin_rom =	37139	;
		9'D197	:	sin_rom =	37305	;
		9'D198	:	sin_rom =	37470	;
		9'D199	:	sin_rom =	37635	;
		9'D200	:	sin_rom =	37800	;
		9'D201	:	sin_rom =	37964	;
		9'D202	:	sin_rom =	38128	;
		9'D203	:	sin_rom =	38292	;
		9'D204	:	sin_rom =	38455	;
		9'D205	:	sin_rom =	38618	;
		9'D206	:	sin_rom =	38781	;
		9'D207	:	sin_rom =	38943	;
		9'D208	:	sin_rom =	39105	;
		9'D209	:	sin_rom =	39266	;
		9'D210	:	sin_rom =	39428	;
		9'D211	:	sin_rom =	39588	;
		9'D212	:	sin_rom =	39749	;
		9'D213	:	sin_rom =	39909	;
		9'D214	:	sin_rom =	40068	;
		9'D215	:	sin_rom =	40227	;
		9'D216	:	sin_rom =	40386	;
		9'D217	:	sin_rom =	40545	;
		9'D218	:	sin_rom =	40703	;
		9'D219	:	sin_rom =	40861	;
		9'D220	:	sin_rom =	41018	;
		9'D221	:	sin_rom =	41175	;
		9'D222	:	sin_rom =	41331	;
		9'D223	:	sin_rom =	41487	;
		9'D224	:	sin_rom =	41643	;
		9'D225	:	sin_rom =	41799	;
		9'D226	:	sin_rom =	41954	;
		9'D227	:	sin_rom =	42108	;
		9'D228	:	sin_rom =	42262	;
		9'D229	:	sin_rom =	42416	;
		9'D230	:	sin_rom =	42569	;
		9'D231	:	sin_rom =	42722	;
		9'D232	:	sin_rom =	42875	;
		9'D233	:	sin_rom =	43027	;
		9'D234	:	sin_rom =	43179	;
		9'D235	:	sin_rom =	43330	;
		9'D236	:	sin_rom =	43481	;
		9'D237	:	sin_rom =	43632	;
		9'D238	:	sin_rom =	43782	;
		9'D239	:	sin_rom =	43931	;
		9'D240	:	sin_rom =	44081	;
		9'D241	:	sin_rom =	44230	;
		9'D242	:	sin_rom =	44378	;
		9'D243	:	sin_rom =	44526	;
		9'D244	:	sin_rom =	44674	;
		9'D245	:	sin_rom =	44821	;
		9'D246	:	sin_rom =	44968	;
		9'D247	:	sin_rom =	45114	;
		9'D248	:	sin_rom =	45260	;
		9'D249	:	sin_rom =	45405	;
		9'D250	:	sin_rom =	45550	;
		9'D251	:	sin_rom =	45695	;
		9'D252	:	sin_rom =	45839	;
		9'D253	:	sin_rom =	45983	;
		9'D254	:	sin_rom =	46126	;
		9'D255	:	sin_rom =	46269	;
		9'D256	:	sin_rom =	46412	;
		9'D257	:	sin_rom =	46554	;
		9'D258	:	sin_rom =	46695	;
		9'D259	:	sin_rom =	46836	;
		9'D260	:	sin_rom =	46977	;
		9'D261	:	sin_rom =	47117	;
		9'D262	:	sin_rom =	47257	;
		9'D263	:	sin_rom =	47396	;
		9'D264	:	sin_rom =	47535	;
		9'D265	:	sin_rom =	47674	;
		9'D266	:	sin_rom =	47812	;
		9'D267	:	sin_rom =	47949	;
		9'D268	:	sin_rom =	48086	;
		9'D269	:	sin_rom =	48223	;
		9'D270	:	sin_rom =	48359	;
		9'D271	:	sin_rom =	48495	;
		9'D272	:	sin_rom =	48630	;
		9'D273	:	sin_rom =	48765	;
		9'D274	:	sin_rom =	48899	;
		9'D275	:	sin_rom =	49033	;
		9'D276	:	sin_rom =	49167	;
		9'D277	:	sin_rom =	49300	;
		9'D278	:	sin_rom =	49432	;
		9'D279	:	sin_rom =	49564	;
		9'D280	:	sin_rom =	49696	;
		9'D281	:	sin_rom =	49827	;
		9'D282	:	sin_rom =	49958	;
		9'D283	:	sin_rom =	50088	;
		9'D284	:	sin_rom =	50217	;
		9'D285	:	sin_rom =	50347	;
		9'D286	:	sin_rom =	50475	;
		9'D287	:	sin_rom =	50604	;
		9'D288	:	sin_rom =	50731	;
		9'D289	:	sin_rom =	50859	;
		9'D290	:	sin_rom =	50985	;
		9'D291	:	sin_rom =	51112	;
		9'D292	:	sin_rom =	51238	;
		9'D293	:	sin_rom =	51363	;
		9'D294	:	sin_rom =	51488	;
		9'D295	:	sin_rom =	51612	;
		9'D296	:	sin_rom =	51736	;
		9'D297	:	sin_rom =	51860	;
		9'D298	:	sin_rom =	51982	;
		9'D299	:	sin_rom =	52105	;
		9'D300	:	sin_rom =	52227	;
		9'D301	:	sin_rom =	52348	;
		9'D302	:	sin_rom =	52469	;
		9'D303	:	sin_rom =	52590	;
		9'D304	:	sin_rom =	52710	;
		9'D305	:	sin_rom =	52829	;
		9'D306	:	sin_rom =	52948	;
		9'D307	:	sin_rom =	53067	;
		9'D308	:	sin_rom =	53185	;
		9'D309	:	sin_rom =	53302	;
		9'D310	:	sin_rom =	53419	;
		9'D311	:	sin_rom =	53535	;
		9'D312	:	sin_rom =	53651	;
		9'D313	:	sin_rom =	53767	;
		9'D314	:	sin_rom =	53882	;
		9'D315	:	sin_rom =	53996	;
		9'D316	:	sin_rom =	54110	;
		9'D317	:	sin_rom =	54223	;
		9'D318	:	sin_rom =	54336	;
		9'D319	:	sin_rom =	54449	;
		9'D320	:	sin_rom =	54561	;
		9'D321	:	sin_rom =	54672	;
		9'D322	:	sin_rom =	54783	;
		9'D323	:	sin_rom =	54893	;
		9'D324	:	sin_rom =	55003	;
		9'D325	:	sin_rom =	55112	;
		9'D326	:	sin_rom =	55221	;
		9'D327	:	sin_rom =	55329	;
		9'D328	:	sin_rom =	55437	;
		9'D329	:	sin_rom =	55544	;
		9'D330	:	sin_rom =	55651	;
		9'D331	:	sin_rom =	55757	;
		9'D332	:	sin_rom =	55862	;
		9'D333	:	sin_rom =	55967	;
		9'D334	:	sin_rom =	56072	;
		9'D335	:	sin_rom =	56176	;
		9'D336	:	sin_rom =	56279	;
		9'D337	:	sin_rom =	56382	;
		9'D338	:	sin_rom =	56485	;
		9'D339	:	sin_rom =	56587	;
		9'D340	:	sin_rom =	56688	;
		9'D341	:	sin_rom =	56789	;
		9'D342	:	sin_rom =	56889	;
		9'D343	:	sin_rom =	56989	;
		9'D344	:	sin_rom =	57088	;
		9'D345	:	sin_rom =	57187	;
		9'D346	:	sin_rom =	57285	;
		9'D347	:	sin_rom =	57382	;
		9'D348	:	sin_rom =	57480	;
		9'D349	:	sin_rom =	57576	;
		9'D350	:	sin_rom =	57672	;
		9'D351	:	sin_rom =	57767	;
		9'D352	:	sin_rom =	57862	;
		9'D353	:	sin_rom =	57957	;
		9'D354	:	sin_rom =	58050	;
		9'D355	:	sin_rom =	58144	;
		9'D356	:	sin_rom =	58236	;
		9'D357	:	sin_rom =	58328	;
		9'D358	:	sin_rom =	58420	;
		9'D359	:	sin_rom =	58511	;
		9'D360	:	sin_rom =	58601	;
		9'D361	:	sin_rom =	58691	;
		9'D362	:	sin_rom =	58781	;
		9'D363	:	sin_rom =	58869	;
		9'D364	:	sin_rom =	58958	;
		9'D365	:	sin_rom =	59045	;
		9'D366	:	sin_rom =	59133	;
		9'D367	:	sin_rom =	59219	;
		9'D368	:	sin_rom =	59305	;
		9'D369	:	sin_rom =	59391	;
		9'D370	:	sin_rom =	59475	;
		9'D371	:	sin_rom =	59560	;
		9'D372	:	sin_rom =	59644	;
		9'D373	:	sin_rom =	59727	;
		9'D374	:	sin_rom =	59809	;
		9'D375	:	sin_rom =	59891	;
		9'D376	:	sin_rom =	59973	;
		9'D377	:	sin_rom =	60054	;
		9'D378	:	sin_rom =	60134	;
		9'D379	:	sin_rom =	60214	;
		9'D380	:	sin_rom =	60293	;
		9'D381	:	sin_rom =	60372	;
		9'D382	:	sin_rom =	60450	;
		9'D383	:	sin_rom =	60528	;
		9'D384	:	sin_rom =	60605	;
		9'D385	:	sin_rom =	60681	;
		9'D386	:	sin_rom =	60757	;
		9'D387	:	sin_rom =	60832	;
		9'D388	:	sin_rom =	60907	;
		9'D389	:	sin_rom =	60981	;
		9'D390	:	sin_rom =	61054	;
		9'D391	:	sin_rom =	61127	;
		9'D392	:	sin_rom =	61199	;
		9'D393	:	sin_rom =	61271	;
		9'D394	:	sin_rom =	61342	;
		9'D395	:	sin_rom =	61413	;
		9'D396	:	sin_rom =	61483	;
		9'D397	:	sin_rom =	61553	;
		9'D398	:	sin_rom =	61621	;
		9'D399	:	sin_rom =	61690	;
		9'D400	:	sin_rom =	61757	;
		9'D401	:	sin_rom =	61824	;
		9'D402	:	sin_rom =	61891	;
		9'D403	:	sin_rom =	61957	;
		9'D404	:	sin_rom =	62022	;
		9'D405	:	sin_rom =	62087	;
		9'D406	:	sin_rom =	62151	;
		9'D407	:	sin_rom =	62215	;
		9'D408	:	sin_rom =	62278	;
		9'D409	:	sin_rom =	62340	;
		9'D410	:	sin_rom =	62402	;
		9'D411	:	sin_rom =	62463	;
		9'D412	:	sin_rom =	62524	;
		9'D413	:	sin_rom =	62584	;
		9'D414	:	sin_rom =	62644	;
		9'D415	:	sin_rom =	62703	;
		9'D416	:	sin_rom =	62761	;
		9'D417	:	sin_rom =	62819	;
		9'D418	:	sin_rom =	62876	;
		9'D419	:	sin_rom =	62932	;
		9'D420	:	sin_rom =	62988	;
		9'D421	:	sin_rom =	63043	;
		9'D422	:	sin_rom =	63098	;
		9'D423	:	sin_rom =	63152	;
		9'D424	:	sin_rom =	63206	;
		9'D425	:	sin_rom =	63259	;
		9'D426	:	sin_rom =	63311	;
		9'D427	:	sin_rom =	63363	;
		9'D428	:	sin_rom =	63414	;
		9'D429	:	sin_rom =	63465	;
		9'D430	:	sin_rom =	63514	;
		9'D431	:	sin_rom =	63564	;
		9'D432	:	sin_rom =	63613	;
		9'D433	:	sin_rom =	63661	;
		9'D434	:	sin_rom =	63708	;
		9'D435	:	sin_rom =	63755	;
		9'D436	:	sin_rom =	63802	;
		9'D437	:	sin_rom =	63847	;
		9'D438	:	sin_rom =	63892	;
		9'D439	:	sin_rom =	63937	;
		9'D440	:	sin_rom =	63981	;
		9'D441	:	sin_rom =	64024	;
		9'D442	:	sin_rom =	64067	;
		9'D443	:	sin_rom =	64109	;
		9'D444	:	sin_rom =	64150	;
		9'D445	:	sin_rom =	64191	;
		9'D446	:	sin_rom =	64232	;
		9'D447	:	sin_rom =	64271	;
		9'D448	:	sin_rom =	64310	;
		9'D449	:	sin_rom =	64349	;
		9'D450	:	sin_rom =	64387	;
		9'D451	:	sin_rom =	64424	;
		9'D452	:	sin_rom =	64461	;
		9'D453	:	sin_rom =	64497	;
		9'D454	:	sin_rom =	64532	;
		9'D455	:	sin_rom =	64567	;
		9'D456	:	sin_rom =	64601	;
		9'D457	:	sin_rom =	64635	;
		9'D458	:	sin_rom =	64668	;
		9'D459	:	sin_rom =	64700	;
		9'D460	:	sin_rom =	64732	;
		9'D461	:	sin_rom =	64763	;
		9'D462	:	sin_rom =	64793	;
		9'D463	:	sin_rom =	64823	;
		9'D464	:	sin_rom =	64853	;
		9'D465	:	sin_rom =	64881	;
		9'D466	:	sin_rom =	64909	;
		9'D467	:	sin_rom =	64937	;
		9'D468	:	sin_rom =	64964	;
		9'D469	:	sin_rom =	64990	;
		9'D470	:	sin_rom =	65016	;
		9'D471	:	sin_rom =	65041	;
		9'D472	:	sin_rom =	65065	;
		9'D473	:	sin_rom =	65089	;
		9'D474	:	sin_rom =	65112	;
		9'D475	:	sin_rom =	65135	;
		9'D476	:	sin_rom =	65157	;
		9'D477	:	sin_rom =	65178	;
		9'D478	:	sin_rom =	65199	;
		9'D479	:	sin_rom =	65219	;
		9'D480	:	sin_rom =	65238	;
		9'D481	:	sin_rom =	65257	;
		9'D482	:	sin_rom =	65275	;
		9'D483	:	sin_rom =	65293	;
		9'D484	:	sin_rom =	65310	;
		9'D485	:	sin_rom =	65326	;
		9'D486	:	sin_rom =	65342	;
		9'D487	:	sin_rom =	65357	;
		9'D488	:	sin_rom =	65372	;
		9'D489	:	sin_rom =	65386	;
		9'D490	:	sin_rom =	65399	;
		9'D491	:	sin_rom =	65412	;
		9'D492	:	sin_rom =	65424	;
		9'D493	:	sin_rom =	65435	;
		9'D494	:	sin_rom =	65446	;
		9'D495	:	sin_rom =	65456	;
		9'D496	:	sin_rom =	65466	;
		9'D497	:	sin_rom =	65475	;
		9'D498	:	sin_rom =	65483	;
		9'D499	:	sin_rom =	65491	;
		9'D500	:	sin_rom =	65498	;
		9'D501	:	sin_rom =	65505	;
		9'D502	:	sin_rom =	65510	;
		9'D503	:	sin_rom =	65516	;
		9'D504	:	sin_rom =	65520	;
		9'D505	:	sin_rom =	65524	;
		9'D506	:	sin_rom =	65528	;
		9'D507	:	sin_rom =	65531	;
		9'D508	:	sin_rom =	65533	;
		9'D509	:	sin_rom =	65534	;
		9'D510	:	sin_rom =	65535	;
		9'D511	:	sin_rom =	65535	;
		default	:	sin_rom =	0	;
		endcase				
	end					
endfunction						
endmodule						
